`ifndef ISA_TYPES_SV
`define ISA_TYPES_SV

typedef enum {
    write_byte,
    write_halfword,
    write_word
} write_width_t;

`endif
