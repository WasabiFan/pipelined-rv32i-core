parameter XLEN = 32;