`ifndef ARCH_CONSTANTS_SV
`define ARCH_CONSTANTS_SV

parameter mem_read_latency = 1'd1;

`endif